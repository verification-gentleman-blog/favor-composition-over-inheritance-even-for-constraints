// Copyright 2018 Tudor Timisescu (verificationgentleman.com)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


package common;

  timeunit 1ns;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "sequence_item.svh"
  `include "sequence_item_stream.svh"

  `include "abstract_test.svh"

  `include "test_all_random.svh"

endpackage
