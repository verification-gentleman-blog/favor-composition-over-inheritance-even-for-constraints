// Copyright 2018 Tudor Timisescu (verificationgentleman.com)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


`include "tests/test_secure_accesses.svh"
`include "tests/test_legal_writes.svh"
`include "tests/test_mapped_addresses.svh"

`include "tests/test_legal_writes_to_mapped_addresses.svh"
`include "tests/test_legal_writes_to_mapped_addresses_in_secure_mode.svh"
