// Copyright 2020 Tudor Timisescu (verificationgentleman.com)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


const bit [31:0] CODE_START_ADDR = 'h0000_0000;
const bit [31:0] CODE_END_ADDR = 'h0fff_ffff;

const bit [31:0] SRAM_START_ADDR = 'h2000_0000;
const bit [31:0] SRAM_END_ADDR = 'h2fff_ffff;

const bit [31:0] PERIPHERAL_START_ADDR = 'h4000_0000;
const bit [31:0] PERIPHERAL_END_ADDR = 'h5fff_ffff;
